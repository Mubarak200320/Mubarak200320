hehbdebheeh
